// vim: set ft=verilog:
`ifndef __CONFIG_H
`define __CONFIG_H

`define MAX_GPIO 7
`define WORD 31

`define LAST_REG 31

`endif
