`include "config.vh"
`include "instructions.vh"

module ram (
  input wire clk,
  input wire en,
  input wire [2:0] write_enable,
  input wire [31:0] addr,
  input wire [31:0] data_in,
  output wire [31:0] data_out
);
  reg [31:0] mem [`RAM_SIZE:0];
  reg [31:0] out;
  integer i;

  wire [31:0] data = mem[addr[12:2]];

  always @(posedge clk) if (en) begin
    out <= addr[1]
      ? (addr[0] ? (data >> 24) : (data >> 16))
      : (addr[0] ? (data >> 8) : data);

    if (write_enable[0]) begin
      mem[addr[12:2]] <= data_in;
    end else if (write_enable[1]) begin
      mem[addr[12:2]] <= addr[1]
        ? {data_in[15:0], data[15:0]}
        : {data[31:16], data_in[15:0]};
    end else if (write_enable[2]) begin
      mem[addr[12:2]] <= addr[1]
        ? (
          addr[0]
          ? {data_in[7:0], data[23:0]}
          : {data[31:24], data[7:0], data[15:0]}
        )
        : (
          addr[0]
          ? {data[31:16], data_in[7:0], data[7:0]}
          : {data[31:8], data_in[7:0]}
        );
    end
  end

  assign data_out = out;
endmodule

module rom (
  input wire clk,
  input wire [31:0] iaddr,
  output wire [31:0] inst
);
  reg [31:0] mem [`ROM_SIZE:0];

  integer i;
  initial $readmemh("firmware/hello.mem", mem);

  assign inst = mem[iaddr >> 2];
endmodule

module iodev (
  input wire clk,
  input wire en,
  input wire [31:0] addr,
  input wire [31:0] data_in,
  output wire [`MAX_GPIO:0] gpio
);
  reg [31:0] gpio_data;

  assign gpio = gpio_data[7:0];

  always @(posedge clk)
    if (en) gpio_data <= data_in;
endmodule

module memory (
  input wire clk,
  input wire [31:0] iaddr,
  input wire [2:0] write_enable,
  input wire [31:0] addr,
  input wire [31:0] data_in,
  output wire [`MAX_GPIO:0] gpio,
  output wire [31:0] data_out,
  output wire [31:0] inst
);
  rom rom (
    .clk(clk),
    .iaddr(iaddr),
    .inst(inst)
  );

  ram ram (
    .clk(clk),
    // ram starts at 0x10000000
    .en(addr[28]),
    .write_enable(write_enable),
    .addr(addr),
    .data_in(data_in),
    .data_out(data_out)
  );

  iodev iodev (
    .clk(clk),
    // iodev starts at 0x20000000
    .en(addr[29]),
    .addr(iaddr),
    .data_in(data_in),
    .gpio(gpio)
  );
endmodule
